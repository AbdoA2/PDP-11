Library ieee;

entity mux2  is  
		port (a, b,s0 : in bit ; x : out bit   );    
	end entity mux2 ;


-- take care of the usage of when else 
architecture  Data_flow of mux2 is
begin
     -- TODO : write the architecture of mux2 
end Data_flow;
